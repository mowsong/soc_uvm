//------------------------------------------------------------
//   Copyright 2010-2012 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------
//
// Class Description:
//
//
class apb_agent_config extends uvm_object;

// UVM Factory Registration Macro
//
`uvm_object_utils(apb_agent_config)

// Virtual Interface
virtual apb_if APB;

//------------------------------------------
// Data Members
//------------------------------------------
// Is the agent active or passive
uvm_active_passive_enum active = UVM_ACTIVE;
// Include the APB functional coverage monitor
bit has_functional_coverage = 0;
// Include the APB RAM based scoreboard
bit has_scoreboard = 0;
//
// Address decode for the select lines:
int no_select_lines = 1;
int apb_index = 0; // Which PSEL is the monitor connected to
bit[31:0] start_address[15:0];
bit[31:0] range[15:0];

bit print_address = 0;

//------------------------------------------
// Methods
//------------------------------------------
// Standard UVM Methods:
extern function new(string name = "apb_agent_config");

extern function string convert2string();

endclass: apb_agent_config

//--------------------------------------------------------------------
//
//--------------------------------------------------------------------
function apb_agent_config::new(string name = "apb_agent_config");
  super.new(name);
endfunction

function string apb_agent_config::convert2string();
  string s;

  s = super.convert2string();
  $sformat(s, "\n");
  $sformat(s, "%s-------------------------------------------------\n", s);
  $sformat(s, "%s  APB AGENT CONFIG                               \n", s);
  $sformat(s, "%s-------------------------------------------------\n", s);
  $sformat(s, "%s  active                  = %s\n", s, active.name());
  $sformat(s, "%s  has_functional_coverage = %b\n", s, has_functional_coverage);
  $sformat(s, "%s  has_scoreboard          = %b\n", s, has_scoreboard);
  if (print_address) begin
  foreach (start_address[i]) begin
    $sformat(s, "%s  start_address[%2d]      = %32h (%32h)\n", 
        s, i, start_address[i], range[i]);
    end
  end
  return s;

endfunction

