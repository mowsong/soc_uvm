package ahb_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "ahb_seq_item.svh"
typedef uvm_sequencer #(ahb_seq_item) ahb_sequencer;
`include "ahb_agent_config.svh"
`include "ahb_driver.svh"
`include "ahb_coverage_monitor.svh"
`include "ahb_monitor.svh"
`include "ahb_agent.svh"

// Utility Sequences

endpackage: ahb_agent_pkg

