module tb_top;
import uvm_pkg::*;

`include "hello_world.svh"

initial begin
  run_test();
end


endmodule

